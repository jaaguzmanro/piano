module piano(wave, t0,t1,t2,t3,t4,t5,t6,t7) 






end module
