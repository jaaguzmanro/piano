module divfreq(freq,chord,clk)

output reg[7:0] freq;
input reg [7:0] chord;
input clk:

    
    
    
    
    
    










endmodule
