module rom(input clk,
                input wire [4:0] addr,
                output reg [3:0] data);


  reg [7:0] rom [0:127];
  always @(negedge clk) begin
    data <= rom[addr];
  end


  initial begin
    rom[0]=00000000;
rom[1]=00000001;
rom[2]=00000010;
rom[3]=00000011;
rom[4]=00000100;
rom[5]=00000101;
rom[6]=00000110;
rom[7]=00000111;
rom[8]=00001000;
rom[9]=00001001;
rom[10]=00001010;
rom[11]=00001011;
rom[12]=00001100;
rom[13]=00001101;
rom[14]=00001110;
rom[15]=00001111;
rom[16]=00010000;
rom[17]=00010001;
rom[18]=00010010;
rom[19]=00010011;
rom[20]=00010100;
rom[21]=00010101;
rom[22]=00010110;
rom[23]=00010111;
rom[24]=00011000;
rom[25]=00011001;
rom[26]=00011010;
rom[27]=00011011;
rom[28]=00011100;
rom[29]=00011101;
rom[30]=00011110;
rom[31]=00011111;
rom[32]=00100000;
rom[33]=00100001;
rom[34]=00100010;
rom[35]=00100011;
rom[36]=00100100;
rom[37]=00100101;
rom[38]=00100110;
rom[39]=00100111;
rom[40]=00101000;
rom[41]=00101001;
rom[42]=00101010;
rom[43]=00101011;
rom[44]=00101100;
rom[45]=00101101;
rom[46]=00101110;
rom[47]=00101111;
rom[48]=00110000;
rom[49]=00110001;
rom[50]=00110010;
rom[51]=00110011;
rom[52]=00110100;
rom[53]=00110101;
rom[54]=00110110;
rom[55]=00110111;
rom[56]=00111000;
rom[57]=00111001;
rom[58]=00111010;
rom[59]=00111011;
rom[60]=00111100;
rom[61]=00111101;
rom[62]=00111110;
rom[63]=00111111;
rom[64]=01000000;
rom[65]=01000001;
rom[66]=01000010;
rom[67]=01000011;
rom[68]=01000100;
rom[69]=01000101;
rom[70]=01000110;
rom[71]=01000111;
rom[72]=01001000;
rom[73]=01001001;
rom[74]=01001010;
rom[75]=01001011;
rom[76]=01001100;
rom[77]=01001101;
rom[78]=01001110;
rom[79]=01001111;
rom[80]=01010000;
rom[81]=01010001;
rom[82]=01010010;
rom[83]=01010011;
rom[84]=01010100;
rom[85]=01010101;
rom[86]=01010110;
rom[87]=01010111;
rom[88]=01011000;
rom[89]=01011001;
rom[90]=01011010;
rom[91]=01011011;
rom[92]=01011100;
rom[93]=01011101;
rom[94]=01011110;
rom[95]=01011111;
rom[96]=01100000;
rom[97]=01100001;
rom[98]=01100010;
rom[99]=01100011;
rom[100]=01100100;
rom[101]=01100101;
rom[102]=01100110;
rom[103]=01100111;
rom[104]=01101000;
rom[105]=01101001;
rom[106]=01101010;
rom[107]=01101011;
rom[108]=01101100;
rom[109]=01101101;
rom[110]=01101110;
rom[111]=01101111;
rom[112]=01110000;
rom[113]=01110001;
rom[114]=01110010;
rom[115]=01110011;
rom[116]=01110100;
rom[117]=01110101;
rom[118]=01110110;
rom[119]=01110111;
rom[120]=01111000;
rom[121]=01111001;
rom[122]=01111010;
rom[123]=01111011;
rom[124]=01111100;
rom[125]=01111101;
rom[126]=01111110;
rom[127]=01111111;
rom[128]=10000000;
rom[129]=10000001;
rom[130]=10000010;
rom[131]=10000011;
rom[132]=10000100;
rom[133]=10000101;
rom[134]=10000110;
rom[135]=10000111;
rom[136]=10001000;
rom[137]=10001001;
rom[138]=10001010;
rom[139]=10001011;
rom[140]=10001100;
rom[141]=10001101;
rom[142]=10001110;
rom[143]=10001111;
rom[144]=10010000;
rom[145]=10010001;
rom[146]=10010010;
rom[147]=10010011;
rom[148]=10010100;
rom[149]=10010101;
rom[150]=10010110;
rom[151]=10010111;
rom[152]=10011000;
rom[153]=10011001;
rom[154]=10011010;
rom[155]=10011011;
rom[156]=10011100;
rom[157]=10011101;
rom[158]=10011110;
rom[159]=10011111;
rom[160]=10100000;
rom[161]=10100001;
rom[162]=10100010;
rom[163]=10100011;
rom[164]=10100100;
rom[165]=10100101;
rom[166]=10100110;
rom[167]=10100111;
rom[168]=10101000;
rom[169]=10101001;
rom[170]=10101010;
rom[171]=10101011;
rom[172]=10101100;
rom[173]=10101101;
rom[174]=10101110;
rom[175]=10101111;
rom[176]=10110000;
rom[177]=10110001;
rom[178]=10110010;
rom[179]=10110011;
rom[180]=10110100;
rom[181]=10110101;
rom[182]=10110110;
rom[183]=10110111;
rom[184]=10111000;
rom[185]=10111001;
rom[186]=10111010;
rom[187]=10111011;
rom[188]=10111100;
rom[189]=10111101;
rom[190]=10111110;
rom[191]=10111111;
rom[192]=11000000;
rom[193]=11000001;
rom[194]=11000010;
rom[195]=11000011;
rom[196]=11000100;
rom[197]=11000101;
rom[198]=11000110;
rom[199]=11000111;
rom[200]=11001000;
rom[201]=11001001;
rom[202]=11001010;
rom[203]=11001011;
rom[204]=11001100;
rom[205]=11001101;
rom[206]=11001110;
rom[207]=11001111;
rom[208]=11010000;
rom[209]=11010001;
rom[210]=11010010;
rom[211]=11010011;
rom[212]=11010100;
rom[213]=11010101;
rom[214]=11010110;
rom[215]=11010111;
rom[216]=11011000;
rom[217]=11011001;
rom[218]=11011010;
rom[219]=11011011;
rom[220]=11011100;
rom[221]=11011101;
rom[222]=11011110;
rom[223]=11011111;
rom[224]=11100000;
rom[225]=11100001;
rom[226]=11100010;
rom[227]=11100011;
rom[228]=11100100;
rom[229]=11100101;
rom[230]=11100110;
rom[231]=11100111;
rom[232]=11101000;
rom[233]=11101001;
rom[234]=11101010;
rom[235]=11101011;
rom[236]=11101100;
rom[237]=11101101;
rom[238]=11101110;
rom[239]=11101111;
rom[240]=11110000;
rom[241]=11110001;
rom[242]=11110010;
rom[243]=11110011;
rom[244]=11110100;
rom[245]=11110101;
rom[246]=11110110;
rom[247]=11110111;
rom[248]=11111000;
rom[249]=11111001;
rom[250]=11111010;
rom[251]=11111011;
rom[252]=11111100;
rom[253]=11111101;
rom[254]=11111110;
rom[255]=11111111;

   end
endmodule
